`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//���������� 4.5 �������� �� HDL ������ minority � ����� �������, a, b, � c,
//� ����� �������, y, ����������� �������� TRUE, ���� �� ����� ���� ������
//����� FALSE.
//////////////////////////////////////////////////////////////////////////////////


module minority(
    input  a, b, c,
    output y
    );
    
    wire [2:0]s ;
    assign s = {a, b, c};
    
    assign y = ((s==3'b000) | (s==3'b001) | (s==3'b010) | (s==3'b100)) ? 1'b1 : 1'b0 ;
     
endmodule
