
// ALU commands
	`define ALU_AND     3'b000
	`define ALU_OR      3'b001
	`define ALU_ADD     3'b010
	`define NOT_USED    3'b011 
	`define ALU_ANDN    3'b100
	`define ALU_ORN		3'b101
	`define ALU_SUB		3'b110
	`define SLT			3'b111
