`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//Упражнение 4.5 Напишите на HDL модуль minority с тремя входами, a, b, и c,
//и одним выходом, y, принимающим значение TRUE, если не менее двух входов
//равны FALSE.
//////////////////////////////////////////////////////////////////////////////////


module minority(
    input  a, b, c,
    output y
    );
    
    wire [2:0]s ;
    assign s = {a, b, c};
    
    assign y = ((s==3'b000) | (s==3'b001) | (s==3'b010) | (s==3'b100)) ? 1'b1 : 1'b0 ;
     
endmodule
